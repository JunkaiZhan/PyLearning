// abd

`define AAAAA hiew.ewew.ewew.ewewewewewe
`define BCG iiuiui.tyty.ytytyty
// `define DJIJ JIJI
`define EEEEE A.b.c.d